-------------------------------------------------------------------------
-- James Gaul
-- CPRE 381
-- Iowa State University
-------------------------------------------------------------------------


-- tb_mux2t1.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file is a testbed for a VDHL 2 to 1 multiplier

--8/31/25 by JAG: Initially Created
-------------------------------------------------------------------------

--Libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.env.all;                -- For hierarchical/external signals
use std.textio.all; 

--Entity Declaration
entity tb_mux2t1 is
  generic(gCLK_HPER   : time := 10 ns);   -- Generic for half of the clock cycle period
end tb_mux2t1;

architecture mixed of tb_mux2t1 is

-- Define the total clock period time
constant cCLK_PER  : time := gCLK_HPER * 2;

--Specifying the component interface
component mux2t1 is
  port(
	i_D0	: in std_logic;
	i_D1	: in std_logic;
	i_S	: in std_logic;
	o_O	: out std_logic);
end component;


-- Create signals for all of the inputs and outputs of the file that you are testing
-- := '0' or := (others => '0') just make all the signals start at an initial value of zero
signal CLK, reset : std_logic := '0';

--input/output signals
signal s_iD0 : std_logic := '0';
signal s_iD1 : std_logic := '0';
signal s_iS : std_logic := '0';
signal s_oO : std_logic;

begin
	DUT0: mux2t1
	port map(
		i_D0	=> s_iD0,
		i_D1	=> s_iD1,
		i_S	=> s_iS,
		o_O	=> s_oO);

  
  --This first process is to setup the clock for the test bench
  P_CLK: process
  begin
    CLK <= '1';         -- clock starts at 1
    wait for gCLK_HPER; -- after half a cycle
    CLK <= '0';         -- clock becomes a 0 (negative edge)
    wait for gCLK_HPER; -- after half a cycle, process begins evaluation again
  end process;


P_TEST_CASES: process
  begin
    wait for gCLK_HPER/2; -- for waveform clarity, I prefer not to change inputs on clk edges

--Case 000
	s_iS	<= '0';	
	s_iD0	<= '0';
	s_iD1	<= '0';
	
	
	wait for gCLK_HPER*2;
	wait for gCLK_HPER*2;

--Case 001
	s_iS	<= '0';
	s_iD0	<= '0';
	s_iD1	<= '1';
	
	wait for gCLK_HPER*2;

--Case 010
	s_iS	<= '0';
	s_iD0	<= '1';
	s_iD1	<= '0';
	
	wait for gCLK_HPER*2;

--Case 011
	s_iS	<= '0';
	s_iD0	<= '1';
	s_iD1	<= '1';
	
	wait for gCLK_HPER*2;

--Case 001
	s_iS	<= '1';
	s_iD0	<= '0';
	s_iD1	<= '0';
	
	wait for gCLK_HPER*2;

--Case 101
	s_iS	<= '1';
	s_iD0	<= '0';
	s_iD1	<= '1';
	
	wait for gCLK_HPER*2;

--Case 110
	s_iS	<= '1';
	s_iD0	<= '1';
	s_iD1	<= '0';
	
	wait for gCLK_HPER*2;

--Case 111
	s_iS	<= '1';
	s_iD0	<= '1';
	s_iD1	<= '1';
	
	wait for gCLK_HPER*2;

wait;
end process;
end mixed;
