Library IEEE;
use IEEE.std_logic_1164.all;

package array32 is
	type array32bits32 is array (0 to 31) of std_logic_vector(31 downto 0);
end package array32;