-------------------------------------------------------------------------
-- James Gaul
-- CPRE 381
-- Iowa State University
-------------------------------------------------------------------------
--Dependencies: RegFile.vhd, addSun_n.vhd, mux2t1_N.vhd
--RISC-V Register system
--Datapath1.vhd
-------------------------------------------------------------------------
--9/24/25 by JAG: Initially Created
-------------------------------------------------------------------------

Library IEEE;
use IEEE.std_logic_1164.all;


entity Datapath2 is
	port(	clock	: in std_logic;
			reset	: in std_logic;
		
			memIn	: in std_logic;
			ALUSrc	: in std_logic; --Determines whether to source from a register(0) or memory/immediate(1)
			--IM_Sw	: in std_logic; --Determines whether to source from immediate (0) or memory(1)

			Imm		: in std_logic_vector(15 downto 0); --16 bit immediate input value

			AddSub	: in std_logic;
			ovflw 	: out std_logic;

		--Register Signals
			Reg_Wr	: in std_logic; --Register write enable
			Rd		: in std_logic_vector(4 downto 0);
			RS1		: in std_logic_vector(4 downto 0);
			RS2		: in std_logic_vector(4 downto 0);

		--Memory Signal
			Mem_Wr	: in std_logic); --Memory write enable
		

end Datapath2;

architecture structural of Datapath2 is
	
   component RegFile is
	port(	clock	: in std_logic;
		reset	: in std_logic;

		RS1Sel	: in std_logic_vector(4 downto 0);
		RS1	: out std_logic_vector(31 downto 0);

		RS2Sel	: in std_logic_vector(4 downto 0);
		RS2	: out std_logic_vector(31 downto 0);

		WrEn	: in std_logic;
		RdSel	: in std_logic_vector(4 downto 0);
		Rd	: in std_logic_vector(31 downto 0));
   end component;

   component addSub_n is
	generic(Comp_Width : integer); -- Generic of type integer for input/output data width.
	port(	nAdd_Sub	: in std_logic;
		i_A		: in std_logic_vector(Comp_Width-1 downto 0);
		i_B		: in std_logic_vector(Comp_Width-1 downto 0);
		o_overflow	: out std_logic;
		o_Sum		: out std_logic_vector(Comp_Width-1 downto 0));
   end component;

   component mux2t1_N is
 	generic(N : integer); -- Generic of type integer for input/output data width. Default value is 32.
 	port(	i_S          : in std_logic;
		i_D0         : in std_logic_vector(N-1 downto 0);
		i_D1         : in std_logic_vector(N-1 downto 0);
		o_O          : out std_logic_vector(N-1 downto 0));
	end component;

component mem is
	generic( 	DATA_WIDTH : natural; 
				ADDR_WIDTH: natural);
	port(	clk		: in std_logic;
			addr 	: in std_logic_vector((ADDR_WIDTH-1) downto 0);
			data 	: in std_logic_vector((DATA_WIDTH-1) downto 0);
			we		: in std_logic := '1';
			q		: out std_logic_vector((DATA_WIDTH -1) downto 0));
end component;
	
component bitExtender16t32 is
	port(	i_sw	: in std_logic;
			i_16bit	: in std_logic_vector(15 downto 0);
			o_32bit	: out std_logic_vector(31 downto 0));
end component;

signal Imm_Ext	: std_logic_vector(31 downto 0)	:= x"00000000";
signal mem_val	: std_logic_vector(31 downto 0)	:= x"00000000";
signal val_in	: std_logic_vector(31 downto 0)	:= x"00000000";

signal sum_b	: std_logic_vector(31 downto 0)	:= x"00000000";

signal Sum_Val	: std_logic_vector(31 downto 0)	:= x"00000000";
signal RS1_Val	: std_logic_vector(31 downto 0)	:= x"00000000";
signal RS2_Val	: std_logic_vector(31 downto 0)	:= x"00000000";
signal RdIn		: std_logic_vector(31 downto 0)	:= x"00000000";

begin
	g_ImmExt: bitExtender16t32
		port map(	i_sw	=> Imm(0),
					i_16bit => Imm,
					o_32bit => Imm_Ext);

	ALUsrcMux:	mux2t1_N
		generic map( N => 32)
		port map(	i_S		=> ALUSrc,
					i_D0	=> RS2_Val,
					i_D1	=> Imm_Ext,
					o_O		=> sum_b);

	RdInMux:	mux2t1_N
		generic map( N => 32)
		port map(	i_S		=> memIn,
					i_D0	=> Sum_Val,
					i_D1	=> mem_val,
					o_O		=> RdIn);

	g_adder: addSub_n
		generic map(	Comp_Width 	=> 32)
		port map(	nAdd_Sub	=> AddSub,
					i_A			=> RS1_Val,
					i_B			=> sum_b,
					o_overflow	=> ovflw,
					o_Sum		=> Sum_Val);

	dmem: mem
		generic map(	DATA_WIDTH	=> 32, 
						ADDR_WIDTH 	=> 10)
		port map(		CLK			=> clock,
						addr		=> Sum_Val(11 downto 2),
						data		=> RS2_Val,
						we			=> Mem_Wr,
						q			=> mem_val);

	g_Reg:	RegFile
		port map(	clock	=> clock,
					reset	=> reset,

					RS1Sel	=> RS1,
					RS1		=> RS1_Val,

					RS2Sel	=> RS2,
					RS2		=> RS2_Val,

					WrEn	=> Reg_Wr,
					RdSel	=> Rd,
					Rd		=> RdIn);
end structural;
