-------------------------------------------------------------------------
-- James Gaul
-- CPRE 381
-- Iowa State University
-------------------------------------------------------------------------


-- tb_mux2t1_N.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbed for an implementation of multiple 2t1 multiplexers

--9/1/25 by JAG: Initially Created
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.env.all;                -- For hierarchical/external signals
use std.textio.all;             -- For basic I/O

-- Usually name your testbench similar to below for clarity tb_<name>
-- TODO: change all instances of tb_TPU_MV_Element to reflect the new testbench.
entity tb_mux2t1_N is
  generic(gCLK_HPER   : time := 10 ns;
          DATA_WIDTH  : integer := 8);   -- Generic for half of the clock cycle period
end tb_mux2t1_N;


architecture mixed of tb_mux2t1_N is

-- Define the total clock period time
constant cCLK_PER  : time := gCLK_HPER * 2;

--Component Interface
component mux2t1_N is
  generic(N : integer); -- Generic of type integer for input/output data width.
  port(i_S          : in std_logic;
       i_D0         : in std_logic_vector(N-1 downto 0);
       i_D1         : in std_logic_vector(N-1 downto 0);
       o_O          : out std_logic_vector(N-1 downto 0));
end component;

--Clock Signal
signal CLK : std_logic := '0';

--Testbed Signals
signal s_iS	: std_logic := '0';
signal s_iD0	: std_logic_vector(DATA_WIDTH-1 downto 0) := x"00";
signal s_iD1	: std_logic_vector(DATA_WIDTH-1 downto 0) := x"00";
signal s_oO	: std_logic_vector(DATA_WIDTH-1 downto 0) := x"00";

begin
	DUT0: mux2t1_N
	generic map (N => DATA_WIDTH)
	port map(
		i_S	=> s_iS,
		i_D0	=> s_iD0,
		i_D1	=> s_iD1,
		o_O	=> s_oO);

--This first process is to setup the clock for the test bench
  P_CLK: process
  begin
    CLK <= '1';         -- clock starts at 1
    wait for gCLK_HPER; -- after half a cycle
    CLK <= '0';         -- clock becomes a 0 (negative edge)
    wait for gCLK_HPER; -- after half a cycle, process begins evaluation again
  end process;

P_TEST_CASES: process
  begin
    wait for gCLK_HPER/2; -- change inputs on clk midpoints

	--Test Case 1:
	s_iS	<= '0';
	s_iD0	<= x"FA";
	s_iD1	<= x"00";
    wait for gCLK_HPER*2;
    

	--Test Case 2:
	s_iS	<= '1';
	s_iD0	<= x"FF";
	s_iD1	<= x"00";
    wait for gCLK_HPER*2;

	--Test Case 2:
	s_iS	<= '0';
	s_iD0	<= x"FF";
	s_iD1	<= x"00";
    wait for gCLK_HPER*2;

	wait;
  end process;
end mixed;