-------------------------------------------------------------------------
-- James Gaul
-- CPRE 381
-- Iowa State University
-------------------------------------------------------------------------


-- onesComp_n.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a ripple carry adder
--9/1/25 by JAG: Initially Created
-------------------------------------------------------------------------

